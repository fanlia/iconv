
module iconv

struct Test {
pub:
	srccode string
	outcode string
	src string
	out string
}

const tests = [
	Test{
		srccode: "UTF8", outcode: "utf-8",
		src: "1111111111111111111111111111111111111111111111111111111111111111" +
			"2222222222222222222222222222222222222222222222222222222222222222" +
			"3333333333333333333333333333333333333333333333333333333333333333" +
			"4444444444444444444444444444444444444444444444444444444444444444" +
			"5555555555555555555555555555555555555555555555555555555555555555" +
			"6666666666666666666666666666666666666666666666666666666666666666" +
			"7777777777777777777777777777777777777777777777777777777777777777" +
			"8888888888888888888888888888888888888888888888888888888888888888" +
			"9999999999999999999999999999999999999999999999999999999999999999" +
			"0000000000000000000000000000000000000000000000000000000000000000",
		out: "1111111111111111111111111111111111111111111111111111111111111111" +
			"2222222222222222222222222222222222222222222222222222222222222222" +
			"3333333333333333333333333333333333333333333333333333333333333333" +
			"4444444444444444444444444444444444444444444444444444444444444444" +
			"5555555555555555555555555555555555555555555555555555555555555555" +
			"6666666666666666666666666666666666666666666666666666666666666666" +
			"7777777777777777777777777777777777777777777777777777777777777777" +
			"8888888888888888888888888888888888888888888888888888888888888888" +
			"9999999999999999999999999999999999999999999999999999999999999999" +
			"0000000000000000000000000000000000000000000000000000000000000000",
	},
	Test{
		srccode: "UTF8", outcode: "utf-8",
		src: "1111111111111111111111111111111111111111111111111111111111111111" +
			"2222222222222222222222222222222222222222222222222222222222222222" +
			"3333333333333333333333333333333333333333333333333333333333333333" +
			"4444444444444444444444444444444444444444444444444444444444444444" +
			"5555555555555555555555555555555555555555555555555555555555555555" +
			"6666666666666666666666666666666666666666666666666666666666666666" +
			"7777777777777777777777777777777777777777777777777777777777777777" +
			"8888888888888888888888888888888888888888888888888888888888888888" +
			"9999999999999999999999999999999999999999999999999999999999999999" +
			"0000000000000000000000000000000000000000000000000000000000000000" +
			"1111111111111111111111111111111111111111111111111111111111111111" +
			"2222222222222222222222222222222222222222222222222222222222222222" +
			"3333333333333333333333333333333333333333333333333333333333333333" +
			"4444444444444444444444444444444444444444444444444444444444444444" +
			"5555555555555555555555555555555555555555555555555555555555555555" +
			"6666666666666666666666666666666666666666666666666666666666666666" +
			"7777777777777777777777777777777777777777777777777777777777777777" +
			"8888888888888888888888888888888888888888888888888888888888888888" +
			"9999999999999999999999999999999999999999999999999999999999999999" +
			"0000000000000000000000000000000000000000000000000000000000000000",
		out: "1111111111111111111111111111111111111111111111111111111111111111" +
			"2222222222222222222222222222222222222222222222222222222222222222" +
			"3333333333333333333333333333333333333333333333333333333333333333" +
			"4444444444444444444444444444444444444444444444444444444444444444" +
			"5555555555555555555555555555555555555555555555555555555555555555" +
			"6666666666666666666666666666666666666666666666666666666666666666" +
			"7777777777777777777777777777777777777777777777777777777777777777" +
			"8888888888888888888888888888888888888888888888888888888888888888" +
			"9999999999999999999999999999999999999999999999999999999999999999" +
			"0000000000000000000000000000000000000000000000000000000000000000" +
			"1111111111111111111111111111111111111111111111111111111111111111" +
			"2222222222222222222222222222222222222222222222222222222222222222" +
			"3333333333333333333333333333333333333333333333333333333333333333" +
			"4444444444444444444444444444444444444444444444444444444444444444" +
			"5555555555555555555555555555555555555555555555555555555555555555" +
			"6666666666666666666666666666666666666666666666666666666666666666" +
			"7777777777777777777777777777777777777777777777777777777777777777" +
			"8888888888888888888888888888888888888888888888888888888888888888" +
			"9999999999999999999999999999999999999999999999999999999999999999" +
			"0000000000000000000000000000000000000000000000000000000000000000",
	},
	Test{
		srccode: "UTF8", outcode: "ISO-8859-1",
		src: "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA" +
			"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA" +
			"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA" +
			"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA" +
			"BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB" +
			"CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC" +
			"dddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddd" +
			"eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee" +
			"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF" +
			"GGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGG" +
			"hhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhh" +
			"iiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiii" +
			"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj" +
			"kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk" +
			"llllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllll" +
			"mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm" +
			"nnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnn" +
			"oooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooo" +
			"pppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppp" +
			"qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq",
		out: "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA" +
			"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA" +
			"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA" +
			"AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA" +
			"BBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBBB" +
			"CCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCCC" +
			"dddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddddd" +
			"eeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeeee" +
			"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF" +
			"GGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGGG" +
			"hhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhhh" +
			"iiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiiii" +
			"jjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjjj" +
			"kkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkkk" +
			"llllllllllllllllllllllllllllllllllllllllllllllllllllllllllllllll" +
			"mmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmmm" +
			"nnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnnn" +
			"oooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooooo" +
			"pppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppppp" +
			"qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq",
	},
]

fn test_iconv() {
	for test in tests {
		cd := iconv.open(test.srccode, test.outcode)
		out := cd.conv_string(test.src)
		assert out == test.out
		cd.close()
	}
}
